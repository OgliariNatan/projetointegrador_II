--INSTITUTO FEDERAL DE SANTA CATARINA

--		PROJETO INTEGRADOR II (2017)

-- 	MENU DE OPÇÃO								RECEBE A SELEÇÃO DE OPÇÃO E DADOS DOS SENSORES
--														EXIBE DADOS NOS DISPLAY 7 SEG	
-- 	AUTORES: 	JEFERSON PEDROSO
--						TARCIS BECHER



LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MENU IS PORT
(
	OPCAO		:	IN	STD_LOGIC_VECTOR (2 DOWNTO 0);
--	DADOS 	:	IN INTEGER;									--AQUI VAI ENTRAR OS DADOS PARA EXIBIR
--	DADOS		: 	IN STD_LOGIC_VECTOR (6 DOWNTO 0);	--DADO PARA TESTE
	DISPLAY0	:	OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
	DISPLAY1	:	OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
	DISPLAY2	:	OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
	DISPLAY3	:	OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
	DISPLAY4	:	OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
	DISPLAY5	:	OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
	DISPLAY6	:	OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
	DISPLAY7	:	OUT STD_LOGIC_VECTOR (6 DOWNTO 0)
);

END MENU;


ARCHITECTURE HARDWARE OF MENU IS 

	BEGIN
	
		WITH OPCAO SELECT
		DISPLAY7		<=		"0001000" WHEN	"001",		--A
								"1000110" WHEN "010",		--C
								"0001100" WHEN "100",		--P
								"1111111" WHEN OTHERS;
								
		WITH OPCAO SELECT
		DISPLAY6		<=		"1000111" WHEN	"001",		--L
								"0100011" WHEN "010",		--o
								"0000100" WHEN "100",		--e
								"1111111" WHEN OTHERS;
								
		WITH OPCAO SELECT
		DISPLAY5		<=		"0000111" WHEN	"001",		--t
								"0101111" WHEN "010",		--r
								"0010010" WHEN "100",		--S
								"1111111" WHEN OTHERS;
								
		WITH OPCAO SELECT
		DISPLAY4		<=		"1100011" WHEN	"001",		--u
								"1111111" WHEN "010",		--'X'
								"0100011" WHEN "100",		--o
								"1111111" WHEN OTHERS;
								

								
								

								
								
		WITH OPCAO SELECT
		DISPLAY1		<=		"0100111" 	WHEN "001",		--c
								--	COR_1	 	WHEN "010",		
							--	"UNID_PESO" WHEN "100",		--g		
								"1111111" 	WHEN OTHERS;			
								
								
		WITH OPCAO SELECT
		DISPLAY0		<=		"0101011" WHEN	"001",		--M
								--COR_0	 WHEN "010",
								--DADOS	 WHEN "010",		
								"0010000" WHEN "100",		--g		
								"1111111" WHEN OTHERS;
								
								
								
								
		
		
	

			
			
END HARDWARE;
		
		
