LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY hc_sr04 IS 
	PORT
	(
	ENABLE	: IN STD_LOGIC;
	ECHO		: IN STD_LOGIC;
	
	TRIGGER	: OUT STD_LOGIC;
	
	);
END hc_sr04;

ARCHITECTURE behavior OF hc_sr04 IS

	BEGIN
	PROCESS()

	END PROCESS;
	
END;