
--		INSTITUTO FEDERAL DE SANTA CATARINA

--		PROJETO INTEGRADOR II (2017)

-- 	DIVISOR DE CLOCK PARA SENSOR HCSR04
--														
-- 	AUTORES: 	JEFERSON	PEDROSO
--						TARCIS	BECHER

--		ABRIL DE 2017

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;




ENTITY cont_pulse IS
	GENERIC (n: POSITIVE := 8);
	PORT(
		CLOCK:		IN STD_LOGIC;
		RST: 			IN STD_LOGIC;
		EN: 			IN STD_LOGIC;
		CONT_PULSE:	OUT STD_LOGIC_VECTOR (n-1 DOWNTO 0)
	);
END cont_pulse;



ARCHITECTURE HARDWARE OF cont_pulse IS

	SIGNAL value: STD_LOGIC_VECTOR(n-1 DOWNTO 0);
	BEGIN
		PROCESS (CLOCK,RST)
		BEGIN
			IF (RST = '1') THEN
				value <= (OTHERS => '0');
			ELSIF (CLOCK'EVENT AND CLOCK='1' AND EN='1') THEN
					value <= value + 1;
			END IF;
		END PROCESS;
		
	CONT_PULSE <= (20-value);
	
END HARDWARE;