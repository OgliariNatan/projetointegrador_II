--INSTITUTO FEDERAL DE SANTA CATARINA

--		PROJETO INTEGRADOR II (2017)

-- 	DECODER 7SEGMENTOS								
--														
-- 	AUTORES: 	JEFERSON PEDROSO
--						TARCIS BECHER

--		ABRIL DE 2017



LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY decode7seg IS PORT
(
	BCD_UNI:		IN	STD_LOGIC_VECTOR (3 DOWNTO 0);
	BCD_DEZ:		IN	STD_LOGIC_VECTOR (3 DOWNTO 0);	
	SEG7_UNI:	OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
	SEG7_DEZ:	OUT STD_LOGIC_VECTOR (6 DOWNTO 0)
);

END decode7seg;


ARCHITECTURE HARDWARE OF decode7seg IS 

	BEGIN
	PROCESS (BCD_UNI)
		BEGIN
		CASE (BCD_UNI) IS
			WHEN "0000" => SEG7_UNI<="1000000";
			WHEN "0001" => SEG7_UNI<="1111001";
			WHEN "0010" => SEG7_UNI<="0100100";
			WHEN "0011" => SEG7_UNI<="0110000";
			WHEN "0100" => SEG7_UNI<="0011001";
			WHEN "0101" => SEG7_UNI<="0010010";
			WHEN "0110" => SEG7_UNI<="0000010";
			WHEN "0111" => SEG7_UNI<="1111000";
			WHEN "1000" => SEG7_UNI<="0000000";
			WHEN "1001" => SEG7_UNI<="0011000";
			WHEN OTHERS	=> SEG7_UNI<="1111111";
		END CASE;		
	END PROCESS;
	
	
	
	
	PROCESS (BCD_DEZ)
		BEGIN
		CASE (BCD_DEZ) IS
			WHEN "0000" => SEG7_DEZ<="1000000";
			WHEN "0001" => SEG7_DEZ<="1111001";
			WHEN "0010" => SEG7_DEZ<="0100100";
			WHEN "0011" => SEG7_DEZ<="0110000";
			WHEN "0100" => SEG7_DEZ<="0011001";
			WHEN "0101" => SEG7_DEZ<="0010010";
			WHEN "0110" => SEG7_DEZ<="0000010";
			WHEN "0111" => SEG7_DEZ<="1111000";
			WHEN "1000" => SEG7_DEZ<="0000000";
			WHEN "1001" => SEG7_DEZ<="0011000";
			WHEN OTHERS	=> SEG7_DEZ<="1111111";
		END CASE;		
	END PROCESS;
	

			
			
END HARDWARE;