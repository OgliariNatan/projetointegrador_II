--INSTITUTO FEDERAL DE SANTA CATARINA

--		PROJETO INTEGRADOR II (2017)

-- 	ENTIDADE MAIN							=>interliga as demais entidades e as conecta ao kit fpga
--														
-- 	AUTORES: 	JEFERSON	PEDROSO
--						TARCIS	BECHER

--		MARÇO DE 2017



LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;



ENTITY MAIN IS PORT
(
	KEY :		IN	STD_LOGIC_VECTOR (3 DOWNTO 0);
	HEX7:	  OUT	STD_LOGIC_VECTOR (6 DOWNTO 0);
	HEX6:	  OUT	STD_LOGIC_VECTOR (6 DOWNTO 0);
	HEX5:	  OUT	STD_LOGIC_VECTOR (6 DOWNTO 0);
	HEX4:	  OUT	STD_LOGIC_VECTOR (6 DOWNTO 0);
	HEX3:	  OUT	STD_LOGIC_VECTOR (6 DOWNTO 0);
	HEX2:	  OUT	STD_LOGIC_VECTOR (6 DOWNTO 0);
	HEX1:	  OUT	STD_LOGIC_VECTOR (6 DOWNTO 0);
	HEX0:	  OUT	STD_LOGIC_VECTOR (6 DOWNTO 0)
);	
	
END MAIN;


ARCHITECTURE HARDWARE OF MAIN IS

	COMPONENT SELETOR						--DECLARAÇÃO DE COMPONENTE (MESMO NOME DA ENTIDADE DE ORIGEM)
		PORT 									--PORT DO COMPONENTE (IGUAL À ENTIDADE DE ORIGEM)
		(
		BOTAO	:	IN	STD_LOGIC;
		SAIDA	: OUT	STD_LOGIC_VECTOR (2 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT MENU
		PORT
		(
		OPCAO		:	IN	STD_LOGIC_VECTOR (2 DOWNTO 0);
--		DADOS 	:	IN INTEGER;									--AQUI VAI ENTRAR OS DADOS PARA EXIBIR
--		DADOS		: 	IN STD_LOGIC_VECTOR (6 DOWNTO 0);	--DADO PARA TESTE
		DISPLAY0	:	OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		DISPLAY1	:	OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		DISPLAY2	:	OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		DISPLAY3	:	OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		DISPLAY4	:	OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		DISPLAY5	:	OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		DISPLAY6	:	OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		DISPLAY7	:	OUT STD_LOGIC_VECTOR (6 DOWNTO 0)
		);
	END COMPONENT;

	
	SIGNAL SEL: STD_LOGIC_VECTOR (2 DOWNTO 0);		--fio para interligar as entidades
	
	
	BEGIN
	
	ROTULO_01:	SELETOR
	
			PORT MAP
			(	KEY(0),
				SEL
			);
				
				
	ROTULO_02: MENU
			
			PORT MAP
			(
			SEL,
	--		DADOS;									--AQUI VAI ENTRAR OS DADOS PARA EXIBIR
			HEX0,
			HEX1,
			HEX2,
			HEX3,
			HEX4,
			HEX5,
			HEX6,
			HEX7
			);
	
	
	
END HARDWARE;