LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;




ENTITY teste_cor IS

	PORT	 ( 
			  );
			  
END teste_cor;




ARCHITECTURE behavior OF teste_cor IS

	

	BEGIN
	
	PROCESS()
	
	
	BEGIN
	
	END PROCESS;
	
END;