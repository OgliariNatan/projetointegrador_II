--INSTITUTO FEDERAL DE SANTA CATARINA

--		PROJETO INTEGRADOR II

-- 	SELETOR DE OPÇÕES

-- 	AUTORES: 	JEFERSON PEDROSO
--						TARCIS BECHER



LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SELETOR IS PORT
(
	BOTAO		:	IN	STD_LOGIC;
	SAIDA		: OUT	STD_LOGIC_VECTOR (2 DOWNTO 0)
);

END SELETOR;


ARCHITECTURE HARDWARE OF SELETOR IS 

	TYPE STATE IS (	CASO_01,				--DECLARAÇÃO DE TIPO
							CASO_02,
							CASO_03);
	
	SIGNAL	ESTADO : STATE; 				--SINAL CHAMADO ESTADO DO TIPO STATE.


	BEGIN	
	
		PROCESSO_SELETOR	:	PROCESS (BOTAO)	--PROCESS CHAMADO PROCESSO_SELETOR SENSIVEL AO BOTAO
			BEGIN
			
			--ESTADO <= CASO_01;				--SETANDO ESTADO INICIAL

			
			IF (BOTAO'EVENT AND BOTAO = '1')	THEN	--QUANDO BOTAO MUDA DE ESTADO AND BOTAO=1
					
				CASE ESTADO IS								--SELEÇÃO DE ESTADOS
					WHEN CASO_01 =>
						ESTADO <= CASO_02;
						
					WHEN CASO_02 =>
						ESTADO <= CASO_03;
						
					WHEN CASO_03 =>
						ESTADO <= CASO_01;
				
				END CASE;
			END IF;
		END PROCESS PROCESSO_SELETOR;
		
		
		WITH ESTADO SELECT							-- CONFIGURA SAIDA DE ACORDO COM O ESTADO
		
			SAIDA <= 	"001" WHEN CASO_01,
							"010" WHEN CASO_02,
							"100" WHEN CASO_03;
--							"000" WHEN OTHERS;
			
			
END HARDWARE;
		
		
